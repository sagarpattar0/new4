module s;
input a;
input b;
input c;

output y;
assign y=a*b
