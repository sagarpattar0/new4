module s;
input a;
input b;
input c;
input d;

output y;
assign y=a*b
