module s;
input a;
input b;
input c;
input d;
input e;

output y;
assign y=a*b
